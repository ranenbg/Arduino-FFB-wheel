CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 75 1918 1031
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
9961490 0
0
2 

2 

0
0
0
24
14 NO PushButton~
191 151 127 0 2 5
0 3 2
0
0 0 4720 0
0
2 B0
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5130 0 0
2
5.90033e-315 5.44746e-315
0
14 NO PushButton~
191 217 127 0 2 5
0 4 2
0
0 0 4720 0
0
2 B1
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
391 0 0
2
5.90033e-315 5.44487e-315
0
14 NO PushButton~
191 353 126 0 2 5
0 6 2
0
0 0 4720 0
0
2 B3
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3124 0 0
2
5.90033e-315 5.44228e-315
0
14 NO PushButton~
191 287 126 0 2 5
0 5 2
0
0 0 4720 0
0
2 B2
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3421 0 0
2
5.90033e-315 5.43969e-315
0
14 NO PushButton~
191 287 181 0 2 5
0 5 9
0
0 0 4720 0
0
2 B6
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8157 0 0
2
5.90033e-315 5.4371e-315
0
14 NO PushButton~
191 353 181 0 2 5
0 6 9
0
0 0 4720 0
0
2 B7
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
5572 0 0
2
5.90033e-315 5.43451e-315
0
14 NO PushButton~
191 217 182 0 2 5
0 4 9
0
0 0 4720 0
0
2 B5
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
8901 0 0
2
5.90033e-315 5.43192e-315
0
14 NO PushButton~
191 151 182 0 2 5
0 3 9
0
0 0 4720 0
0
2 B4
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
7361 0 0
2
5.90033e-315 5.42933e-315
0
14 NO PushButton~
191 152 289 0 2 5
0 3 7
0
0 0 4720 0
0
3 B12
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4747 0 0
2
5.90033e-315 5.42414e-315
0
14 NO PushButton~
191 218 289 0 2 5
0 4 7
0
0 0 4720 0
0
3 B13
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
972 0 0
2
5.90033e-315 5.41896e-315
0
14 NO PushButton~
191 354 288 0 2 5
0 6 7
0
0 0 4720 0
0
3 B15
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3472 0 0
2
5.90033e-315 5.41378e-315
0
14 NO PushButton~
191 288 288 0 2 5
0 5 7
0
0 0 4720 0
0
3 B14
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
9998 0 0
2
5.90033e-315 5.4086e-315
0
14 NO PushButton~
191 288 233 0 2 5
0 5 8
0
0 0 4720 0
0
3 B10
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3536 0 0
2
5.90033e-315 5.40342e-315
0
14 NO PushButton~
191 354 233 0 2 5
0 6 8
0
0 0 4720 0
0
3 B11
-10 -20 11 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4597 0 0
2
5.90033e-315 5.39824e-315
0
14 NO PushButton~
191 218 234 0 2 5
0 4 8
0
0 0 4720 0
0
2 B9
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3835 0 0
2
5.90033e-315 5.39306e-315
0
14 NO PushButton~
191 152 234 0 2 5
0 3 8
0
0 0 4720 0
0
2 B8
-7 -20 7 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3670 0 0
2
5.90033e-315 5.38788e-315
0
11 Terminal:A~
194 87 152 0 1 3
0 2
0
0 0 49648 0
2 D6
-23 -4 -9 4
2 J1
-7 -23 7 -15
0
3 D6;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
5616 0 0
2
5.90033e-315 5.37752e-315
0
11 Terminal:A~
194 176 81 0 1 3
0 3
0
0 0 49648 270
2 D4
-7 -17 7 -9
2 J5
-7 -23 7 -15
0
3 D4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
9323 0 0
2
5.90033e-315 5.36716e-315
0
11 Terminal:A~
194 243 81 0 1 3
0 4
0
0 0 49648 270
2 A4
-7 -17 7 -9
2 J6
-7 -23 7 -15
0
3 A4;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
317 0 0
2
5.90033e-315 5.3568e-315
0
11 Terminal:A~
194 313 81 0 1 3
0 5
0
0 0 49648 270
2 A5
-6 -17 8 -9
2 J7
-7 -23 7 -15
0
3 A5;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
3108 0 0
2
5.90033e-315 5.34643e-315
0
11 Terminal:A~
194 382 81 0 1 3
0 6
0
0 0 49648 270
3 D12
-10 -17 11 -9
2 J8
-7 -23 7 -15
0
4 D12;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
4299 0 0
2
5.90033e-315 5.32571e-315
0
11 Terminal:A~
194 87 313 0 1 3
0 7
0
0 0 49648 0
2 D5
-23 -4 -9 4
2 J4
-7 -23 7 -15
0
3 D5;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
9672 0 0
2
5.90033e-315 5.30499e-315
0
11 Terminal:A~
194 87 260 0 1 3
0 8
0
0 0 49648 0
2 D8
-23 -4 -9 4
2 J3
-7 -23 7 -15
0
3 D8;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
7876 0 0
2
5.90033e-315 5.26354e-315
0
11 Terminal:A~
194 87 207 0 1 3
0 9
0
0 0 49648 0
2 D7
-23 -4 -9 4
2 J2
-7 -23 7 -15
0
3 D7;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 J
6369 0 0
2
5.90033e-315 0
0
32
2 0 7 0 0 8192 0 9 0 0 4 3
135 297
125 297
125 313
2 0 7 0 0 0 0 10 0 0 4 3
201 297
192 297
192 313
2 0 7 0 0 8192 0 12 0 0 4 3
271 296
263 296
263 313
1 2 7 0 0 4224 0 22 11 0 0 4
93 313
330 313
330 296
337 296
2 0 8 0 0 8192 0 16 0 0 8 3
135 242
125 242
125 260
2 0 8 0 0 0 0 15 0 0 8 3
201 242
192 242
192 260
2 0 8 0 0 8192 0 13 0 0 8 3
271 241
263 241
263 260
1 2 8 0 0 4224 0 23 14 0 0 4
93 260
330 260
330 241
337 241
2 0 9 0 0 8192 0 8 0 0 12 3
134 190
125 190
125 207
2 0 9 0 0 0 0 7 0 0 12 3
200 190
192 190
192 207
2 0 9 0 0 8192 0 5 0 0 12 3
270 189
263 189
263 207
1 2 9 0 0 4224 0 24 6 0 0 4
93 207
330 207
330 189
336 189
2 0 2 0 0 8192 0 4 0 0 16 3
270 134
263 134
263 152
2 0 2 0 0 0 0 2 0 0 16 3
200 135
192 135
192 152
2 0 2 0 0 0 0 1 0 0 16 3
134 135
125 135
125 152
2 1 2 0 0 12416 0 3 17 0 0 4
336 134
330 134
330 152
93 152
1 0 6 0 0 4096 0 3 0 0 20 2
370 134
382 134
1 0 6 0 0 0 0 6 0 0 20 2
370 189
382 189
1 0 6 0 0 0 0 14 0 0 20 2
371 241
382 241
1 1 6 0 0 4224 0 21 11 0 0 3
382 87
382 296
371 296
1 0 5 0 0 4096 0 4 0 0 24 2
304 134
313 134
1 0 5 0 0 0 0 5 0 0 24 2
304 189
313 189
1 0 5 0 0 0 0 13 0 0 24 2
305 241
313 241
1 1 5 0 0 4224 0 20 12 0 0 3
313 87
313 296
305 296
1 0 4 0 0 4096 0 2 0 0 28 2
234 135
243 135
1 0 4 0 0 0 0 7 0 0 28 2
234 190
243 190
1 0 4 0 0 0 0 15 0 0 28 2
235 242
243 242
1 1 4 0 0 4224 0 19 10 0 0 3
243 87
243 297
235 297
1 0 3 0 0 4096 0 1 0 0 32 2
168 135
176 135
1 0 3 0 0 0 0 8 0 0 32 2
168 190
176 190
1 0 3 0 0 0 0 16 0 0 32 2
169 242
176 242
1 1 3 0 0 4224 0 18 9 0 0 3
176 87
176 297
169 297
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
